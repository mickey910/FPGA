library verilog;
use verilog.vl_types.all;
entity noblocking_vlg_vec_tst is
end noblocking_vlg_vec_tst;
