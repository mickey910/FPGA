library verilog;
use verilog.vl_types.all;
entity blocking_vlg_vec_tst is
end blocking_vlg_vec_tst;
