library verilog;
use verilog.vl_types.all;
entity part3_vlg_vec_tst is
end part3_vlg_vec_tst;
