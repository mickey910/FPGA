library verilog;
use verilog.vl_types.all;
entity ip_counter_vlg_vec_tst is
end ip_counter_vlg_vec_tst;
